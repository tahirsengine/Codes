// megafunction wizard: %LPM_MULT%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_mult 

// ============================================================
// File Name: mult1.v
// Megafunction Name(s):
// 			lpm_mult
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 18.0.0 Build 614 04/24/2018 SJ Lite Edition
// ************************************************************

//Copyright (C) 2018  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details.

module mult1 (
	dataa,
	datab,
	result);

	input	[1:0]  dataa;
	input	[1:0]  datab;
	output	[4:0]  result;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: AutoSizeResult NUMERIC "0"
// Retrieval info: PRIVATE: B_isConstant NUMERIC "0"
// Retrieval info: PRIVATE: ConstantB NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX 10"
// Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "0"
// Retrieval info: PRIVATE: Latency NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: SignedMult NUMERIC "0"
// Retrieval info: PRIVATE: USE_MULT NUMERIC "1"
// Retrieval info: PRIVATE: ValidConstant NUMERIC "0"
// Retrieval info: PRIVATE: WidthA NUMERIC "2"
// Retrieval info: PRIVATE: WidthB NUMERIC "2"
// Retrieval info: PRIVATE: WidthP NUMERIC "5"
// Retrieval info: PRIVATE: aclr NUMERIC "0"
// Retrieval info: PRIVATE: clken NUMERIC "0"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: PRIVATE: optimize NUMERIC "0"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_HINT STRING "DEDICATED_MULTIPLIER_CIRCUITRY=YES,MAXIMIZE_SPEED=5"
// Retrieval info: CONSTANT: LPM_REPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MULT"
// Retrieval info: CONSTANT: LPM_WIDTHA NUMERIC "2"
// Retrieval info: CONSTANT: LPM_WIDTHB NUMERIC "2"
// Retrieval info: CONSTANT: LPM_WIDTHP NUMERIC "5"
// Retrieval info: USED_PORT: dataa 0 0 2 0 INPUT NODEFVAL "dataa[1..0]"
// Retrieval info: USED_PORT: datab 0 0 2 0 INPUT NODEFVAL "datab[1..0]"
// Retrieval info: USED_PORT: result 0 0 5 0 OUTPUT NODEFVAL "result[4..0]"
// Retrieval info: CONNECT: @dataa 0 0 2 0 dataa 0 0 2 0
// Retrieval info: CONNECT: @datab 0 0 2 0 datab 0 0 2 0
// Retrieval info: CONNECT: result 0 0 5 0 @result 0 0 5 0
// Retrieval info: GEN_FILE: TYPE_NORMAL mult1.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult1.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult1.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult1.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult1_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult1_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
